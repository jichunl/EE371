// The 4-bit ripple down counter

`include "DFilpFlop.v"

module ripple_down_counter 
	(input 	wire		clk_i 
	,input 	wire		reset_i
	,output reg	[3:0] 	q_o
	);

	wire q0, q1, q2, q3;
	
	
	
	
endmodule

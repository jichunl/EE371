// This is the module that controls the pressure (ie. fill and evacuate the 
//	chamber) inside the interlock
// Input:
//	clk_i: the clock that this module runs on
//	rst_i: the signal that resets this module
// 	
// Output:
//	fill_o: the signal 
// 	evac_o:
